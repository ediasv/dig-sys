library ieee;
use ieee.std_logic_1164.all;

entity cont_999 is
  port (
    i_clk : in std_logic;
    o_clk : out std_logic
  );
end entity;

architecture behavioral of cont_999 is
  signal internal_clk : std_logic;
begin
end architecture behavioral;
