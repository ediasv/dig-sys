library ieee;
use ieee.std_logic_1164.all;

entity lab4 is 
  port();
end entity;
