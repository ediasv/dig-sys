library ieee;
use ieee.std_logic_1164.all;

entity eduardo is
  port (
    :w;w
  );
end entity eduardo;

architecture rtl of eduardo is
begin
end architecture rtl;
